oscconf_inst : oscconf PORT MAP (
		oscena	 => oscena_sig,
		osc	 => osc_sig
	);
